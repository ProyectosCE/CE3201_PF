 module Instruction_Memory(
 
 input logic [31:0] a,
 
 output logic [31:0] rd
 
 );
 
 
endmodule 

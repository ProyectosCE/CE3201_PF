module Gambling_Tec(




);



endmodule

module marioSprite(input [9:0] pixel_x,
						 input [9:0] pixel_y,
						 input [9:0] posx,
						 input [9:0] posy,
						 output logic [23:0] RGB,
						 output visible);
			

logic [23:0] RGB_i, RGB_ii;

logic [3:0]  sprite_i [0:31] [0:31]   = 
'{'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b0011, 4'b1101, 4'b1101, 4'b0101, 4'b0111, 4'b1101, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1101, 4'b1101, 4'b1100, 4'b0101, 4'b1000, 4'b0111, 4'b1100, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1101, 4'b1100, 4'b1100, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1101, 4'b1100, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1100, 4'b1100, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1100, 4'b0011, 4'b0001, 4'b0001, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b0010, 4'b0010, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b1110, 4'b1110, 4'b0010, 4'b0001, 4'b0100, 4'b0001, 4'b0010, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b1110, 4'b0001, 4'b0100, 4'b0001, 4'b0001, 4'b1110, 4'b0100, 4'b0010, 4'b0001, 4'b0100, 4'b0001, 4'b0010, 4'b0100, 4'b0110, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b1110, 4'b0001, 4'b1110, 4'b0001, 4'b0001, 4'b0001, 4'b0100, 4'b0100, 4'b1110, 4'b1110, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0110, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b1110, 4'b1110, 4'b1110, 4'b0001, 4'b0100, 4'b0100, 4'b0001, 4'b0110, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b0110, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0001, 4'b1110, 4'b1110, 4'b1110, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0110, 4'b1110, 4'b1110, 4'b0100, 4'b0100, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b0011, 4'b0001, 4'b0101, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b0101, 4'b0101, 4'b0101, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1100, 4'b1100, 4'b1100, 4'b1100, 4'b1100, 4'b1100, 4'b0011, 4'b0011, 4'b0101, 4'b0101, 4'b0101, 4'b0010, 4'b0101, 4'b0010, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1100, 4'b1101, 4'b1101, 4'b1101, 4'b1101, 4'b1010, 4'b1010, 4'b1101, 4'b1101, 4'b1010, 4'b0000, 4'b0101, 4'b0010, 4'b0010, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1100, 4'b0101, 4'b0101, 4'b0101, 4'b1100, 4'b1100, 4'b1001, 4'b1001, 4'b1100, 4'b1100, 4'b1001, 4'b0101, 4'b0010, 4'b0010, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b0101, 4'b0010, 4'b0010, 4'b0101, 4'b0101, 4'b0011, 4'b0011, 4'b1011, 4'b1011, 4'b0011, 4'b0011, 4'b1011, 4'b0101, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0010, 4'b0010, 4'b0010, 4'b0010, 4'b0010, 4'b0101, 4'b1011, 4'b1000, 4'b1000, 4'b1011, 4'b1011, 4'b1000, 4'b1010, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0010, 4'b0010, 4'b0010, 4'b0010, 4'b0010, 4'b0101, 4'b1011, 4'b1000, 4'b1000, 4'b1011, 4'b1011, 4'b1010, 4'b0101, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0010, 4'b0010, 4'b0010, 4'b0101, 4'b1011, 4'b1011, 4'b1011, 4'b1011, 4'b1011, 4'b1010, 4'b0101, 4'b1000, 4'b0101, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0101, 4'b0101, 4'b0101, 4'b1001, 4'b1001, 4'b1011, 4'b1011, 4'b1011, 4'b1010, 4'b0101, 4'b0101, 4'b0101, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0101, 4'b0101, 4'b1010, 4'b1010, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1010, 4'b0101, 4'b0101, 4'b0101, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0101, 4'b0101, 4'b1010, 4'b1010, 4'b1010, 4'b1010, 4'b1010, 4'b1010, 4'b1010, 4'b1010, 4'b0101, 4'b0101, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0101, 4'b1000, 4'b0101, 4'b0101, 4'b1010, 4'b1010, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0101, 4'b0101, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}};


logic [3:0] RGB_i_encoded_i;

assign RGB_i_encoded_i = sprite_i [pixel_y-posy][pixel_x-posx];

//color table
always_comb
	case(RGB_i_encoded_i)
	4'h0: RGB_i = 24'h464646;
	4'h1: RGB_i = 24'h000000;
	4'h2: RGB_i = 24'hFFFFFF;
	4'h3: RGB_i = 24'h00007b;
	4'h4: RGB_i = 24'ha8d9ff;
	4'h5: RGB_i = 24'h134e6a;
	4'h6: RGB_i = 24'h005882;
	4'h7: RGB_i = 24'h15abb0;
	4'h8: RGB_i = 24'h59e6ea;
	4'h9: RGB_i = 24'hc58452;
	4'hA: RGB_i = 24'h964602;
	4'hB: RGB_i = 24'hffc28f;
	4'hC: RGB_i = 24'h1700c9;
	4'hD: RGB_i = 24'h4B36FF;
	4'hE: RGB_i = 24'h7d73ff;
	default:  RGB_i = 24'h464646;
	endcase

	
logic n_back_i;
assign n_back_i = (RGB_i_encoded_i == 4'b0000);	
logic visible_i;
assign visible_i = (~n_back_i & posx[0]) & ((pixel_x >=  posx) & (pixel_x < posx + 10'd32)) & (( pixel_y >=  posy) & (pixel_y < posy + 10'd32));	




logic [3:0]  sprite [0:31] [0:31]   = 
'{'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b0011, 4'b1101, 4'b1101, 4'b1111, 4'b0111, 4'b1101, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1101, 4'b1101, 4'b1100, 4'b1111, 4'b1000, 4'b0111, 4'b1100, 4'b0011, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1101, 4'b1100, 4'b1100, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1101, 4'b1100, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1100, 4'b1100, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1100, 4'b0011, 4'b0001, 4'b0001, 4'b1110, 4'b0010, 4'b0010, 4'b1110, 4'b0010, 4'b0010, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0011, 4'b0001, 4'b0001, 4'b1110, 4'b1110, 4'b0010, 4'b0001, 4'b0100, 4'b0001, 4'b0010, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b1110, 4'b0001, 4'b0100, 4'b0001, 4'b0001, 4'b1110, 4'b0100, 4'b0010, 4'b0001, 4'b0100, 4'b0001, 4'b0010, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b1110, 4'b0001, 4'b1110, 4'b0001, 4'b0001, 4'b0001, 4'b0100, 4'b0100, 4'b1110, 4'b1110, 4'b0100, 4'b0100, 4'b0100, 4'b0100, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b1110, 4'b1110, 4'b1110, 4'b0001, 4'b0100, 4'b0100, 4'b0001, 4'b0101, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0001, 4'b1110, 4'b1110, 4'b1110, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0101, 4'b1110, 4'b1110, 4'b0100, 4'b0100, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b1110, 4'b0101, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b1100, 4'b1100, 4'b0011, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1101, 4'b1101, 4'b0011, 4'b1100, 4'b1111, 4'b0010, 4'b0010, 4'b1111, 4'b1111, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1100, 4'b1101, 4'b1101, 4'b1101, 4'b1111, 4'b0010, 4'b0010, 4'b0010, 4'b0010, 4'b0010, 4'b1111, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0011, 4'b1100, 4'b1100, 4'b1101, 4'b1101, 4'b1111, 4'b0010, 4'b1111, 4'b0010, 4'b0010, 4'b1111, 4'b1111, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b1010, 4'b0011, 4'b1100, 4'b1100, 4'b1101, 4'b1101, 4'b1111, 4'b0010, 4'b0010, 4'b1111, 4'b1111, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b1010, 4'b1010, 4'b0011, 4'b1100, 4'b1100, 4'b0011, 4'b0011, 4'b1111, 4'b1111, 4'b1111, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b1010, 4'b1001, 4'b1010, 4'b0011, 4'b0011, 4'b0011, 4'b1000, 4'b1000, 4'b1011, 4'b1000, 4'b1010, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b1010, 4'b1001, 4'b1011, 4'b1011, 4'b1011, 4'b1011, 4'b1011, 4'b1011, 4'b1011, 4'b1001, 4'b1010, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b1010, 4'b1001, 4'b1011, 4'b1011, 4'b1011, 4'b1011, 4'b1010, 4'b1001, 4'b1010, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b1010, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1001, 4'b1010, 4'b1001, 4'b1010, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b1010, 4'b1010, 4'b1010, 4'b1010, 4'b1010, 4'b1010, 4'b1010, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0101, 4'b0101, 4'b0101, 4'b0101, 4'b0101, 4'b0001, 4'b0101, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0101, 4'b0101, 4'b0101, 4'b0101, 4'b1000, 4'b0001, 4'b1000, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0001, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}, 
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000},
'{4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000, 4'b0000}};


logic [3:0] RGB_encoded;

assign RGB_encoded = sprite [pixel_y-posy][pixel_x-posx];

//color table
always_comb
	case(RGB_encoded)
	4'h0: RGB_ii = 24'h464646;
	4'h1: RGB_ii = 24'h000000;
	4'h2: RGB_ii = 24'hFFFFFF;
	4'h3: RGB_ii = 24'h00007b;
	4'h4: RGB_ii = 24'ha8d9ff;
	4'h5: RGB_ii = 24'h134e6a;
	4'h6: RGB_ii = 24'h005882;
	4'h7: RGB_ii = 24'h15abb0;
	4'h8: RGB_ii = 24'h59e6ea;
	4'h9: RGB_ii = 24'hc58452;
	4'hA: RGB_ii= 24'h964602;
	4'hB: RGB_ii = 24'hffc28f;
	4'hC: RGB_ii = 24'h1700c9;
	4'hD: RGB_ii = 24'h4B36FF;
	4'hE: RGB_ii = 24'h7d73ff;
	4'hF: RGB_ii = 24'h046777;
	default:  RGB_ii = 24'h464646;
	endcase

	
logic n_back;
assign n_back = (RGB_encoded == 4'b0000);	
logic visible_ii;
assign visible_ii = (~n_back & ~posx[0]) & ((pixel_x >=  posx) & (pixel_x < posx + 10'd32)) & (( pixel_y >=  posy) & (pixel_y < posy + 10'd32));	


assign visible = visible_i | visible_ii;

assign RGB = posx[0] ? RGB_i: RGB_ii;


endmodule

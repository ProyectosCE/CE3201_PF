module Bit_cell(



);


endmodule 
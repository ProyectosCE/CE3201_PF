module Deslizador(


);


endmodule

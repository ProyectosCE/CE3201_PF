module Rom_tile (
	input  logic [9:0] Q_X, Q_Y,
	output logic visible,
	output logic [7:0] R, G, B
);

logic [2:0] sprite_i [0:14][0:31] = '{
    '{3'b000, 3'b001, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000},
    '{3'b000, 3'b000, 3'b001, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000},
    '{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
    '{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b000, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001},
    '{3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b001, 3'b000, 3'b000, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000},
    '{3'b001, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b010, 3'b010, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000},
    '{3'b000, 3'b001, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b001},
    '{3'b000, 3'b000, 3'b000, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b001, 3'b000, 3'b001, 3'b000, 3'b000, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b000, 3'b000, 3'b001, 3'b001, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000},
    '{3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b001, 3'b000, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010},
    '{3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010},
    '{3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010},
    '{3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b010, 3'b000, 3'b001, 3'b001, 3'b000, 3'b001, 3'b001, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010},
    '{3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010},
    '{3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b001, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010},
    '{3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010}
};

logic [4:0] local_x;
logic [3:0] local_y;
logic [2:0] pixel;

assign local_x = Q_X % 32;
assign local_y = Q_Y % 15;
assign pixel = sprite_i[local_y][local_x];

// Define el área donde se debe ver el sprite
logic Area_div;
assign Area_div = ((Q_X > 420 && Q_X < 440) || (Q_X > 520 && Q_X < 540)) &&
                  (Q_Y > 160 && Q_Y < 460);

// RGB con color solo si estamos dentro del área
always_comb begin
	if (Area_div) begin
		case (pixel)
			3'b001: begin R = 8'hFF; G = 8'hFF; B = 8'h00; end // amarillo
			3'b010: begin R = 8'h00; G = 8'h00; B = 8'hFF; end // azul
			default: begin R = 8'h00; G = 8'h00; B = 8'h00; end // negro
		endcase
	end else begin
		R = 8'h00; G = 8'h00; B = 8'h00; // fondo fuera del área
	end
end

assign visible = Area_div;

endmodule
